module cpu(input wire clk, reset);
//Procesador sin memoria de datos de un solo ciclo


endmodule
